/*
 *  TOPPERS/ASP Kernel
 *      Toyohashi Open Platform for Embedded Real-Time Systems/
 *      Advanced Standard Profile Kernel
 * 
 *  Copyright (C) 2015 by Ushio Laboratory
 *              Graduate School of Engineering Science, Osaka Univ., JAPAN
 *  Copyright (C) 2015,2016 by Embedded and Real-Time Systems Laboratory
 *              Graduate School of Information Science, Nagoya Univ., JAPAN
 * 
 *  上記著作権者は，以下の(1)〜(4)の条件を満たす場合に限り，本ソフトウェ
 *  ア（本ソフトウェアを改変したものを含む．以下同じ）を使用・複製・改
 *  変・再配布（以下，利用と呼ぶ）することを無償で許諾する．
 *  (1) 本ソフトウェアをソースコードの形で利用する場合には，上記の著作
 *      権表示，この利用条件および下記の無保証規定が，そのままの形でソー
 *      スコード中に含まれていること．
 *  (2) 本ソフトウェアを，ライブラリ形式など，他のソフトウェア開発に使
 *      用できる形で再配布する場合には，再配布に伴うドキュメント（利用
 *      者マニュアルなど）に，上記の著作権表示，この利用条件および下記
 *      の無保証規定を掲載すること．
 *  (3) 本ソフトウェアを，機器に組み込むなど，他のソフトウェア開発に使
 *      用できない形で再配布する場合には，次のいずれかの条件を満たすこ
 *      と．
 *    (a) 再配布に伴うドキュメント（利用者マニュアルなど）に，上記の著
 *        作権表示，この利用条件および下記の無保証規定を掲載すること．
 *    (b) 再配布の形態を，別に定める方法によって，TOPPERSプロジェクトに
 *        報告すること．
 *  (4) 本ソフトウェアの利用により直接的または間接的に生じるいかなる損
 *      害からも，上記著作権者およびTOPPERSプロジェクトを免責すること．
 *      また，本ソフトウェアのユーザまたはエンドユーザからのいかなる理
 *      由に基づく請求からも，上記著作権者およびTOPPERSプロジェクトを
 *      免責すること．
 * 
 *  本ソフトウェアは，無保証で提供されているものである．上記著作権者お
 *  よびTOPPERSプロジェクトは，本ソフトウェアに関して，特定の使用目的
 *  に対する適合性も含めて，いかなる保証も行わない．また，本ソフトウェ
 *  アの利用により直接的または間接的に生じたいかなる損害に関しても，そ
 *  の責任を負わない．
 * 
 *  $Id: tSIOPortTarget.cdl 1799 2023-04-01 00:50:30Z ertl-komori $
 */

/*
 * シリアルインタフェースドライバのターゲット依存部
 * のコンポーネント記述
 */

/*
 * ボードに関する定義
 */
import_C("frdm_mcxn947.h");
import_C("MCXNx4x.h");

/*
 * USART用 簡易SIOドライバ
 */
import("tUsart.cdl");

/*
 * シリアルインタフェースドライバのターゲット依存部の本体（シリアルイ
 * ンタフェースドライバとSIOドライバを接続する部分）のセルタイプ
 */
celltype tSIOPortTargetMain {
    /*
     *  シリアルインタフェースドライバとの結合
     */
    [inline]   entry    sSIOPort    eSIOPort;
    [optional] call     siSIOCBR    ciSIOCBR;

    /*
     *  SIOドライバとの結合
     */
    call              sSIOPort    cSIOPort;
    [inline] entry    siSIOCBR    eiSIOCBR;

    /*
     *  割込み要求ライン操作のための結合
     */
    call    sInterruptRequest    cInterruptRequest;
};

/*
 * シリアルインタフェースドライバのターゲット依存部（複合コンポーネン
 * ト）のセルタイプ
 */
[active]
composite tSIOPortTarget {
    /*
     * シリアルインタフェースドライバとの結合
     */
    entry              sSIOPort    eSIOPort;
    [optional] call    siSIOCBR    ciSIOCBR;

    /*
     * 属性の定義
     */
    attr {
        uintptr_t baseAddress;            /* ベースアドレス */
        uintptr_t flexcommAddress;        /* Flexcommアドレス */
        uint32_t  index;                  /* USARTインデックス */
        INTNO     interruptNumber;        /* 割込み番号 */
        PRI       isrPriority = 1;        /* ISR優先度 */
        PRI       interruptPriority = -2; /* 割込み優先度 */
    };

    /*
     * SIOドライバ
     */
    cell tUsart Usart {
        baseAddress     = composite.baseAddress;
        flexcommAddress = composite.flexcommAddress;
        index           = composite.index;
        ciSIOCBR        = SIOPortMain.eiSIOCBR;
    };

    /*
     * シリアルインタフェースドライバのターゲット依存部の本体
     */
    cell tSIOPortTargetMain SIOPortMain {
        ciSIOCBR          => composite.ciSIOCBR;
        cSIOPort          = Usart.eSIOPort;
        cInterruptRequest = InterruptRequest.eInterruptRequest;
    };
    composite.eSIOPort => SIOPortMain.eSIOPort;

    /*
     * SIOの割込みサービスルーチンと割込み要求ライン
     */
    cell tISR ISRInstance {
        interruptNumber = composite.interruptNumber;
        isrPriority     = composite.isrPriority;
        ciISRBody       = Usart.eiISR;
    };
    cell tInterruptRequest InterruptRequest {
        interruptNumber   = composite.interruptNumber;
        interruptPriority = composite.interruptPriority;
    };
};

/*
 * シリアルインタフェースドライバのターゲット依存部のプロトタイプ
 */
[prototype]
cell tSIOPortTarget SIOPortTarget1 {
    baseAddress     = C_EXP("MCXNx4x_LPUART4_BASE");
    flexcommAddress = C_EXP("MCXNx4x_LP_FLEXCOMM4_BASE");
    index           = C_EXP("4");
    interruptNumber = C_EXP("MCXNx4x_LP_FLEXCOMM4_IRQ + 16");
};

/* 
[prototype]
cell tSIOPortTarget SIOPortTarget2 {
    baseAddress     = C_EXP("MCXNx4x_LPUART1_BASE");
    flexcommAddress = C_EXP("MCXNx4x_LP_FLEXCOMM1_BASE");
    index           = C_EXP("1");
    interruptNumber = C_EXP("MCXNx4x_LP_FLEXCOMM1_IRQ + 16");
};

[prototype]
cell tSIOPortTarget SIOPortTarget3 {
    baseAddress     = C_EXP("MCXNx4x_LPUART2_BASE");
    flexcommAddress = C_EXP("MCXNx4x_LP_FLEXCOMM2_BASE");
    index           = C_EXP("2");
    interruptNumber = C_EXP("MCXNx4x_LP_FLEXCOMM2_IRQ + 16");
};

[prototype]
cell tSIOPortTarget SIOPortTarget4 {
    baseAddress     = C_EXP("MCXNx4x_LPUART3_BASE");
    flexcommAddress = C_EXP("MCXNx4x_LP_FLEXCOMM3_BASE");
    index           = C_EXP("3");
    interruptNumber = C_EXP("MCXNx4x_LP_FLEXCOMM3_IRQ + 16");
};

[prototype]
cell tSIOPortTarget SIOPortTarget5 {
    baseAddress     = C_EXP("MCXNx4x_LPUART4_BASE");
    flexcommAddress = C_EXP("MCXNx4x_LP_FLEXCOMM4_BASE");
    index           = C_EXP("4");
    interruptNumber = C_EXP("MCXNx4x_LP_FLEXCOMM4_IRQ + 16");
};

[prototype]
cell tSIOPortTarget SIOPortTarget6 {
    baseAddress     = C_EXP("MCXNx4x_LPUART5_BASE");
    flexcommAddress = C_EXP("MCXNx4x_LP_FLEXCOMM5_BASE");
    index           = C_EXP("5");
    interruptNumber = C_EXP("MCXNx4x_LP_FLEXCOMM5_IRQ + 16");
};

[prototype]
cell tSIOPortTarget SIOPortTarget7 {
    baseAddress     = C_EXP("MCXNx4x_LPUART6_BASE");
    flexcommAddress = C_EXP("MCXNx4x_LP_FLEXCOMM6_BASE");
    index           = C_EXP("6");
    interruptNumber = C_EXP("MCXNx4x_LP_FLEXCOMM6_IRQ + 16");
};

[prototype]
cell tSIOPortTarget SIOPortTarget8 {
    baseAddress     = C_EXP("MCXNx4x_LPUART7_BASE");
    flexcommAddress = C_EXP("MCXNx4x_LP_FLEXCOMM7_BASE");
    index           = C_EXP("7");
    interruptNumber = C_EXP("MCXNx4x_LP_FLEXCOMM7_IRQ + 16");
};
*/
